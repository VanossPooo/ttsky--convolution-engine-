module convolution_engine (
	input  wire [7:0] ui_in,    // Number to be put in matrix
    	output wire [7:0] uo_out,   // Dedicated outputs
    	input  wire [7:0] uio_in,   // Size
    	output wire [7:0] uio_out,  // IOs: Output path
    	output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    	input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    	input  wire       clk,      // clock
    	input  wire       rst_n );    // reset_n - low to reset


Buffer U1 ();
Padding U2 ();

endmodule